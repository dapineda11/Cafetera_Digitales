library verilog;
use verilog.vl_types.all;
entity Expreso_vlg_vec_tst is
end Expreso_vlg_vec_tst;
